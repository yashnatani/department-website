CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 110 10 100 9
0 74 1024 471
7 5.000 V
7 5.000 V
3 GND
50 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 74 1024 471
144179219 0
0
6 Title:
5 Name:
0
0
0
16
7 Ground~
168 438 304 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
11 Signal Gen~
195 482 141 0 64 64
0 7 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1112014847 0 1077936128
1015598705 814313567 814313567 981668463 1017370379 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162691
20
0 50 0 3 0.0167 1e-009 1e-009 0.001 0.02 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/3V
-15 -30 13 -22
2 V4
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(0 3 16.7m 1n 1n 1m 20m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
11 Signal Gen~
195 386 143 0 64 64
0 8 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1112014847 0 1077936128
1008971033 814313567 814313567 981668463 1017370379 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162722
20
0 50 0 3 0.00999 1e-009 1e-009 0.001 0.02 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/3V
-15 -30 13 -22
2 V8
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(0 3 9.99m 1n 1n 1m 20m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
11 Signal Gen~
195 295 148 0 64 64
0 9 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1112014847 0 1077936128
995769377 814313567 814313567 981668463 1017370379 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162720
20
0 50 0 3 0.00333 1e-009 1e-009 0.001 0.02 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/3V
-15 -30 13 -22
2 V9
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(0 3 3.33m 1n 1n 1m 20m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
4 SCR~
219 527 223 0 3 7
0 4 7 3
0
0 0 848 180
6 2N6241
-53 0 -11 8
4 SCR3
-46 -10 -18 -2
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-126
7

0 2 3 1 2 3 1 0
88 0 0 256 1 0 0 0
3 SCR
5394 0 0
0
0
4 SCR~
219 445 222 0 3 7
0 5 8 3
0
0 0 848 180
6 2N6241
-53 0 -11 8
4 SCR2
-46 -10 -18 -2
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-126
7

0 2 3 1 2 3 1 0
88 0 0 256 1 0 0 0
3 SCR
7734 0 0
0
0
4 SCR~
219 371 221 0 3 7
0 6 9 3
0
0 0 848 180
6 2N6241
-53 0 -11 8
4 SCR1
-46 -10 -18 -2
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-126
7

0 2 3 1 2 3 1 0
88 0 0 256 1 1 0 0
3 SCR
9914 0 0
0
0
6 Diode~
219 519 264 0 2 5
0 2 4
0
0 0 848 90
6 1N5406
8 0 50 8
2 D3
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
6 DO-201
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3747 0 0
0
0
6 Diode~
219 438 264 0 2 5
0 2 5
0
0 0 848 90
6 1N5406
8 0 50 8
2 D2
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
6 DO-201
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3549 0 0
0
0
6 Diode~
219 364 263 0 2 5
0 2 6
0
0 0 848 90
6 1N5406
8 0 50 8
2 D1
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
6 DO-201
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7931 0 0
0
0
7 Ground~
168 165 370 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
11 Signal Gen~
195 124 489 0 20 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1120403456
1012557331
20
1 50 0 100 0.01333 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 90
9 -100/100V
27 3 90 11
2 V3
52 -7 66 1
0
0
43 %D %1 %2 DC 0 SIN(0 100 50 13.33m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
11 Signal Gen~
195 209 428 0 20 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1120403456
1004170870
20
1 50 0 100 0.006666 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 90
9 -100/100V
27 3 90 11
2 V2
52 -7 66 1
0
0
43 %D %1 %2 DC 0 SIN(0 100 50 6.666m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3834 0 0
0
0
11 Signal Gen~
195 51 396 0 19 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1120403456
20
1 50 0 100 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 90
9 -100/100V
27 3 90 11
2 V1
52 -7 66 1
0
0
38 %D %1 %2 DC 0 SIN(0 100 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
9 Resistor~
219 717 170 0 2 5
0 3 10
0
0 0 880 0
3 100
-10 -12 11 -4
2 R5
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 812 239 0 3 5
0 2 10 -1
0
0 0 880 90
3 500
4 -1 25 7
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
23
3 1 3 0 0 8320 0 5 15 0 0 3
519 211
519 170
699 170
0 1 2 0 0 4096 0 0 1 19 0 2
438 282
438 298
1 0 4 0 0 8320 0 12 0 0 16 3
127 456
127 249
519 249
1 2 5 0 0 8320 0 13 9 0 0 4
212 395
212 246
438 246
438 254
1 0 6 0 0 8320 0 14 0 0 18 3
54 363
54 248
364 248
1 2 2 0 0 12288 0 11 13 0 0 4
165 364
165 256
222 256
222 395
1 2 2 0 0 0 0 11 12 0 0 4
165 364
165 360
137 360
137 456
1 2 2 0 0 0 0 11 14 0 0 4
165 364
165 360
64 360
64 363
1 2 7 0 0 8320 0 2 5 0 0 4
513 136
542 136
542 217
532 217
1 2 8 0 0 8320 0 3 6 0 0 6
417 138
453 138
453 206
457 206
457 216
450 216
1 2 9 0 0 8320 0 4 7 0 0 6
326 143
353 143
353 238
386 238
386 215
376 215
1 1 2 0 0 8320 0 8 16 0 0 4
519 274
519 278
812 278
812 257
2 1 2 0 0 0 0 4 11 0 0 5
326 153
330 153
330 356
165 356
165 364
2 2 2 0 0 0 0 3 2 0 0 6
417 148
453 148
453 167
521 167
521 146
513 146
2 2 2 0 0 0 0 4 3 0 0 6
326 153
357 153
357 169
425 169
425 148
417 148
1 2 4 0 0 0 0 5 8 0 0 2
519 235
519 254
1 2 5 0 0 0 0 6 9 0 0 4
437 234
437 246
438 246
438 254
1 2 6 0 0 0 0 7 10 0 0 4
363 233
363 245
364 245
364 253
1 1 2 0 0 0 0 9 8 0 0 4
438 274
438 282
519 282
519 274
1 1 2 0 0 0 0 10 9 0 0 4
364 273
364 282
438 282
438 274
3 3 3 0 0 0 0 6 5 0 0 4
437 210
437 203
519 203
519 211
3 3 3 0 0 0 0 7 6 0 0 4
363 209
363 202
437 202
437 210
2 2 10 0 0 4224 0 15 16 0 0 3
735 170
812 170
812 221
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0.02 0.1 0.001 0.001
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
3605398 8550464 100 100 0 0
77 66 977 246
0 406 1024 738
974 66
77 66
977 66
977 246
0 0
0.0997335 0.0200422 120 -120 0.0799578 0.0799578
12401 0
4 0.03 1e+009
8
699 170
0 3 0 0 2	0 1 0 0
532 217
0 7 0 0 3	0 9 0 0
452 216
0 8 0 0 5	0 10 0 0
363 233
0 6 0 0 1	0 18 0 0
437 235
0 5 0 0 1	0 17 0 0
519 235
0 4 0 0 1	0 16 0 0
812 221
0 10 0 0 2	0 23 0 0
376 215
0 9 0 0 5	0 11 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
