CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
0 74 1024 406
8  5.000 V
8  5.000 V
3 GND
50 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 74 1024 406
144179219 0
0
6 Title:
5 Name:
0
0
0
20
10 Polar Cap~
219 758 187 0 2 5
0 4 3
0
0 0 848 270
3 1uF
10 4 31 12
2 C1
14 -6 28 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8953 0 0
0
0
9 Inductor~
219 139 140 0 2 5
0 11 8
0
0 0 848 0
5 0.1mH
-18 -17 17 -9
2 L3
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
9 Inductor~
219 139 109 0 2 5
0 12 9
0
0 0 848 0
5 0.1mH
-18 -17 17 -9
2 L2
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
9 Inductor~
219 138 81 0 2 5
0 13 10
0
0 0 848 0
5 0.1mH
-18 -17 17 -9
2 L4
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
7 Ground~
168 129 315 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
11 Signal Gen~
195 222 222 0 20 64
0 11 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
1012557331
20
1 50 0 250 0.01333 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V3
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 SIN(0 250 50 13.33m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
11 Signal Gen~
195 131 222 0 20 64
0 12 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
1004157985
20
1 50 0 250 0.00666 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V2
-7 -40 7 -32
0
0
42 %D %1 %2 DC 0 SIN(0 250 50 6.66m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
11 Signal Gen~
195 45 222 0 19 64
0 13 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
20
1 50 0 250 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 250 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
9 Inductor~
219 641 120 0 2 5
0 15 14
0
0 0 848 0
5 0.5mH
-18 -17 17 -9
2 L1
-7 -27 7 -19
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
6 Diode~
219 456 245 0 2 5
0 3 6
0
0 0 848 90
5 DIODE
11 0 46 8
2 D6
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
7931 0 0
0
0
6 Diode~
219 542 139 0 2 5
0 5 15
0
0 0 848 90
5 DIODE
11 0 46 8
2 D5
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
9325 0 0
0
0
6 Diode~
219 371 247 0 2 5
0 3 7
0
0 0 848 90
5 DIODE
11 0 46 8
2 D4
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
8903 0 0
0
0
6 Diode~
219 443 140 0 2 5
0 6 15
0
0 0 848 90
5 DIODE
11 0 46 8
2 D3
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3834 0 0
0
0
6 Diode~
219 506 249 0 2 5
0 3 5
0
0 0 848 90
5 DIODE
11 0 46 8
2 D2
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3363 0 0
0
0
6 Diode~
219 356 142 0 2 5
0 7 15
0
0 0 848 90
5 DIODE
11 0 46 8
2 D1
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
7668 0 0
0
0
9 Resistor~
219 189 139 0 2 5
0 8 5
0
0 0 880 0
2 1m
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 189 108 0 2 5
0 9 6
0
0 0 880 0
2 1m
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 188 80 0 2 5
0 10 7
0
0 0 880 0
2 1m
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 802 187 0 2 5
0 3 4
0
0 0 880 90
4 16.5
1 0 29 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 707 118 0 2 5
0 14 4
0
0 0 880 0
2 2M
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 1 0 0
1 R
4871 0 0
0
0
25
2 1 3 0 0 8192 0 1 19 0 0 4
757 194
757 213
802 213
802 205
0 1 4 0 0 12288 0 0 1 16 0 4
728 118
728 110
757 110
757 177
2 0 5 0 0 12416 0 16 0 0 23 4
207 139
344 139
344 165
542 165
2 0 6 0 0 4224 0 17 0 0 24 4
207 108
430 108
430 165
443 165
2 0 7 0 0 4224 0 18 0 0 25 4
206 80
343 80
343 156
356 156
2 1 8 0 0 12416 0 2 16 0 0 4
157 140
163 140
163 139
171 139
2 1 9 0 0 12416 0 3 17 0 0 4
157 109
163 109
163 108
171 108
2 1 10 0 0 12416 0 4 18 0 0 4
156 81
162 81
162 80
170 80
1 1 11 0 0 12416 0 6 2 0 0 6
253 217
257 217
257 148
113 148
113 140
121 140
1 1 12 0 0 8320 0 7 3 0 0 6
162 217
166 217
166 114
113 114
113 109
121 109
1 1 13 0 0 8320 0 8 4 0 0 4
76 217
102 217
102 81
120 81
1 2 2 0 0 8320 0 5 6 0 0 5
129 309
129 247
261 247
261 227
253 227
1 2 2 0 0 0 0 5 7 0 0 5
129 309
129 247
170 247
170 227
162 227
2 1 2 0 0 0 0 8 5 0 0 5
76 227
102 227
102 301
129 301
129 309
0 1 3 0 0 4224 0 0 19 19 0 3
456 265
802 265
802 205
2 2 4 0 0 4224 0 20 19 0 0 3
725 118
802 118
802 169
2 1 14 0 0 4224 0 9 20 0 0 4
659 120
681 120
681 118
689 118
0 1 15 0 0 4224 0 0 9 21 0 4
443 121
615 121
615 120
623 120
1 1 3 0 0 0 0 10 14 0 0 4
456 255
456 267
506 267
506 259
1 1 3 0 0 0 0 12 10 0 0 4
371 257
371 263
456 263
456 255
2 2 15 0 0 0 0 13 11 0 0 4
443 130
443 121
542 121
542 129
2 2 15 0 0 0 0 15 13 0 0 4
356 132
356 122
443 122
443 130
1 2 5 0 0 0 0 11 14 0 0 4
542 149
542 231
506 231
506 239
1 2 6 0 0 0 0 13 10 0 0 4
443 150
443 227
456 227
456 235
1 2 7 0 0 0 0 15 12 0 0 4
356 152
356 229
371 229
371 237
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0.02 0.1 0.002 0.002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
6685644 1079360 100 100 0 0
77 66 977 186
0 74 161 144
977 66
77 66
977 66
977 186
0 0
0.5 0 270 -270 0.5 540
12385 0
4 0.01 10000
0
6685668 8550976 100 100 0 0
77 66 977 246
0 406 1024 738
977 66
77 66
977 66
977 180
0 0
0.080621 0.020621 300 -80 0.079379 0.079379
12409 0
2 0.01 100
4
764 118
0 4 0 0 1	0 16 0 0
356 156
0 7 0 0 3	0 5 0 0
443 153
0 6 0 0 1	0 24 0 0
542 152
0 5 0 0 1	0 23 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
