CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 74 1024 582
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 74 1024 582
144441362 0
0
6 Title:
5 Name:
0
0
0
7
7 Ground~
168 235 429 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
11 Signal Gen~
195 140 347 0 20 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
1012557331
20
1 50 0 250 0.01333 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V3
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 SIN(0 250 50 13.33m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
11 Signal Gen~
195 140 277 0 20 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
1004170870
20
1 50 0 250 0.006666 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V2
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 SIN(0 250 50 6.666m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
11 Signal Gen~
195 139 207 0 19 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
20
1 50 0 250 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 250 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
9 Resistor~
219 486 200 0 4 5
0 3 2 0 -1
0
0 0 880 0
4 100k
-14 -14 14 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 393 201 0 4 5
0 4 2 0 -1
0
0 0 880 0
4 100k
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
9 Resistor~
219 305 201 0 4 5
0 5 2 0 -1
0
0 0 880 0
4 100k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
9
2 1 2 0 0 12416 0 5 1 0 0 5
504 200
508 200
508 415
235 415
235 423
1 1 3 0 0 4224 0 2 5 0 0 4
171 342
460 342
460 200
468 200
2 0 2 0 0 128 0 6 0 0 5 4
411 201
415 201
415 418
235 418
1 1 4 0 0 4224 0 3 6 0 0 4
171 272
367 272
367 201
375 201
2 1 2 0 0 128 0 7 1 0 0 5
323 201
327 201
327 415
235 415
235 423
1 1 5 0 0 4224 0 4 7 0 0 4
170 202
279 202
279 201
287 201
2 2 2 0 0 0 0 3 4 0 0 4
171 282
178 282
178 212
170 212
2 2 2 0 0 0 0 2 3 0 0 4
171 352
179 352
179 282
171 282
2 1 2 0 0 128 0 2 1 0 0 3
171 352
235 352
235 423
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.5 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
4916172 8546880 100 100 0 0
77 66 977 186
0 478 1024 738
114 66
77 66
977 66
977 126
0 0
0.00493333 0 300 0 0.5 0.5
12409 0
2 0.02 100
3
172 272
0 4 0 0 1	0 4 0 0
191 202
0 5 0 0 1	0 6 0 0
173 342
0 3 0 0 1	0 2 0 0
3867596 8550976 100 100 0 0
77 66 977 246
0 406 1024 738
977 66
77 66
977 66
977 246
0 0
0.005 0 300 0 0.005 0.005
12409 0
4 0.001 100
1
239 202
0 3 0 0 1	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
